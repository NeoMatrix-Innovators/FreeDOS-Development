Begin3
Language:    SV, 850
Title:       switchar
Description: Visa och s�tt DOS switchar
Keywords:    freedos
End
