FD-REPOv1	Build time: 1645361091	Ljudverktyg	5
adplay	1.6b	musikseplare f�r flera format som anv�nder OPL2/3-ljud	1197d98e
cdp	A4 (rev A)	Audio CD-spelare f�r DOS kommandorad	76265c51
dosmid	0.9.5a	MIDI-spelare f�r m�nga synthesizrar (AWE, MPU-401, OPL...)	a4ba39bd
mplayer	1.0rc2 (rev A)	MPlayer �r en videospelare porterad fr�n Linux.	79c7bf85
opencp	2.6.0pre6 (rev A)	OpenCubic Player �r en musikspelare f�r m�nga format (mp3,wav,mid...)	fb37a44c
