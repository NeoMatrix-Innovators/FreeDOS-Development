Begin3
Language:    SV, 850
Title:       PCISLEEP
Description: PCISLEEP listar och s�ver pci-kort.
Keywords:    PCISleep, pci, card, vga, sova, lista
End
