Begin3
Language:    SV, 850
Title:       UDVD2
Description: CD/DVD UltraDMA-enhetsdrivrutin
Keywords:    cd, disk, dma, drivrutin, dvd, ultra
End
