Begin3
Language:    SV, 850
Title:       Biew
Description: Biew �r en bin�r/hexadecimal visare/redigerare. (kr�ver i686+)
Keywords:    Biew, bin�r, hexadecimal, visare, redigerarer
End
