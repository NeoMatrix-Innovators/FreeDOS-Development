Begin3
Language:    SV, 850
Title:       Testdisk (och Photorec)
Description: Testdisk kontrollerar partitioner/startsektorer p� diskar; Photorec �terst�ller m�nga typer av data
Keywords:    testdisk, photorec, data, �terst�ll, test
End
