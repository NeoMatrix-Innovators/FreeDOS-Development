Begin3
Language:    SV, 850
Title:       Doszip Commander
Description: En liten LFN-medveten filhanterare med inbyggd zip-uppackare. Den �r byggd med JWasm och OpenWatcom. Inkluderar fullst�ndig k�llkod f�r DOS och Windows
Keywords:    DOS FreeDOS
End
