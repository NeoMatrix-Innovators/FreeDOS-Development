Begin3
Language:    SV, 850
Title:       UnZip
Description: Ett fildekomprimeringsverktyg i stil med PKUNZIP.
Keywords:    freedos, unzip, infozip, pkunzip
End
