Begin3
Language:    SV, 850
Title:       DISKCOMP
Description: Diskj�mf�reelseverktyg
Keywords:    diskcomp, j�mf�r, diskar
End
