Begin3
Language:    SV, 850
Title:       GNU chcp
Description: LOADFONT (GNUCHCP) �ndrar EGA-/VGA-bitmappstypsnitt p� sk�rmen i textl�ge.
Keywords:    loadfont gnuchcp bitmapp typsnitt ega vga sk�rm
End
