Begin3
Language:    SV, 850
Title:       SHSUCDX
Description: En fri CDROM-extender f�r DOS
Keywords:    mscdex, shsucdex, fdcdex, cdrom, atapicdd, xcdrom
End
