Begin3
Language:    SV, 850
Title:       Search
Description: Hittar filer p� din dator
Keywords:    freedos, s�k
End
