Begin3
Language:    SV, 850
Title:       GNU bc
Description: bc �r ett numerisk behandlingsspr�k med godtycklig precision. Syntaxen liknar C, men skiljer sig p� ett flertal omr�den. Det har st�d f�r interaktiv k�rning av satser. bc�r ett verktyg som inkluderas i standardutkastet POSIX P1003.2/D11.
Keywords:    kalkylator, bc, gnubc
End
