Begin3
Language:    SV, 850
Title:       COMP
Description: J�mf�r filer och visa deras skillnader
Keywords:    j�mf�r, comp, filj�mf�relse
End
