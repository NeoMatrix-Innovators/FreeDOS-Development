Begin3
Language:    SV, 850
Title:       Gopherus
Description: En fri, (16-bitars) konsolll�gesklient f�r gopher f�r flera plattformar
Summary:     Gopherus �r en fri gopher-klient f�r konsoll�ge f�r flera plattformar s� som DOS, LInux och Windows. Den tillhandah�ller ett klassiskt textgr�nssnitt till gopher-rymden. �ven om den i f�rsta hand �r riktad mot DOS finns porteringar ocks� f�r Windows och Linux. Dessa anv�nder SDL2 f�r att emulera en pseudo-terminal. (16-bitarsversion)
Keywords:    gopher n�tverk n�tverk
End
