Begin3
Language:    SV, 850
Title:       MSEDIT
Description: Mateusz Saucy Editor
Keywords:    textredigerare
End
