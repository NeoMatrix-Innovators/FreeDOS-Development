Begin3
Language:    SV, 850
Title:       aefdisk
Description: Kommandoradsdrivet diskpartitioneringsverktyg f�r DOS (portat f�r Open Watcom)
Keywords:    dos fdisk partition
End
