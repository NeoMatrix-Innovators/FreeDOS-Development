Begin3
Language:    SV, 850
Title:       Dillo
Description: En grafisk webbl�sare k�nd f�r sin hastighet och lilla minnesavtryck.
Keywords:    dillo, webb, www, l�sare
End
