FD-REPOv1	Build time: 1645361091	Unix-liknande verktyg	16
cal	1.07a	Kalenderprogram, i stil med UNIX cal	25b7be9c
du	1.0a	Visa diskanv�ndning, i stil med du under UNIX	b7833017
gnubc	1.02a	bc �r ett numerisk behandlingsspr�k med godtycklig precision. Syntaxen liknar C, men skiljer sig p� ett flertal omr�den. Det har st�d f�r interaktiv k�rning av satser. bc�r ett verktyg som inkluderas i standardutkastet POSIX P1003.2/D11.	be361cdb
gnused	4.2.2a	GNU sed �r en GNU-implementation av POSIX str�mredigerarer `sed'.	f8b2f576
grep	2.0a	grep genoms�ker filer (eller standard in) efter rader som matcar ett givet m�nster. M�nstret kan vara ett regulj�rt uttryck eller en bokstavlig str�ng.	1831fda3
head	1.0a	Visar en del av en fil	c10358ad
less	291a	Less �r ett program i stil med more, men vilket l�ter dig g� bak�t i filen s� v�l som fram�t. Less m�ste heller inte l�sa hela indatafilen innan den startar, s� f�r st�rre indatafiler startar det upp snabbare �n textredigerare som vi.	6536b9c0
md5sum	3.0a	Ber�knar MD5 kontrollsummor	71586e3c
nro	1.2a	En textbehandlare i stil med nroff i UNIX	b9ece9dd
sleep	1.0a	sleep liknar UNIX-verktyget med samma namn. sleep kan anv�ndas f�r att pausa k�rningen av kommandofiler en studn. sleep ger tillbaka tid till operativsystem som har st�d f�r det. sleep k�nner igen och respekterar DOS switchar.	f1322eee
tee	2.0.3a	Sparar en kopia av dess indata till en fil, medan en kopia skrivs ut p� stdout	dc1ecfcf
touch	1.4.4a	S�tter datum- och tidst�mplar p� filer likt touch i *nix	b4fc87a3
trch	3.1g	�vers�tter tecken. Detta kan anv�ndas med programmet UNIX2DOS, men kan �vers�tta fler tecken. [Liknar, men �r inte samma som, tr i UNIX.] (inkluderar Cats GNU LGPL)	4b117090
uptimec	2.60a	Rapporterar k�rtid, �ven inuti DOSEmu. Liknar uptime i UNIX.	55e9c9c4
which	2.1a	which �r ett verktyg fr�n UNIX-v�rlden som l�ter anv�ndare hitta k�rbara filer i katalogerna listade i milj�variabeln PATH. Fullt st�d f�r jokertecken, relativa s�kv�gare, valfria fildetaljer (storlek, datum). Anv�ndardefinierbara program�ndelser, kodsides-korreka tids-/datumformatering. Nytt DOS sitchar-st�d.	0a9c224b
xgrep	1.03a	Snabb UNIX-liknande `grep'-klon med st�d f�r regulj�ra uttryck	6801a74d
