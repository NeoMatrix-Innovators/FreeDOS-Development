Begin3
Language:    SV, 850
Title:       DOG
Description: Ett alternativs command.com-skal, i stil med FreeCOM, men annorlunda.
Keywords:    kommando, skal
End
