Begin3
Language:    SV, 850
Title:       CTMouse
Description: FreeDOS musdrivrutin
Keywords:    Mus, hjul
End
