Begin3
Language:    SV, 850
Title:       SRDISK (resizeable RAM disk)
Description: Ramdisk som kan �ndra storlek. Srdisk �r en snabb och kan anv�nd mer �n 32MB XMS och EMS-minne. Storleken p� disket kan �ndras utan att starta och eller att f�rlora inneh�ll. Kompatibel med diskcopy.
Keywords:    ut�kning, verktyg, ramdisk
End
