Begin3
Language:    SV, 850
Title:       WhichFAT
Description: K�rnst�d f�r FAT32 identifiering och FAT-typdetektering (12-32) per enhet
Keywords:    freedos, fat, disk
End
