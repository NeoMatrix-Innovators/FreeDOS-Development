Begin3
Language:    SV, 850
Title:       xkeyb
Description: Tangentbordsdrivrutin f�r internationellt st�d. Inkluderar ocks� KEYMAN + KLIB + LISTXDEF + SCANKBD
Keywords:    keyb, tangentbord, drivrutin
End
