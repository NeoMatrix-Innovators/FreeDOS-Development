Begin3
Language:    SV, 850
Title:       Floppy Bird
Description: Floppy Bird �r en klon av det �k�nda Flappy Bird skriven i 16 -bitars (x86) assembler. Med andra or fungerar det p� RENT KISEL och kr�ver inte ett underliggande operativsystem, det �r ett operativsystem i sig.
Keywords:    spel, action
End
