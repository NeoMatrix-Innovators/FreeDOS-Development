Begin3
Language:    SV, 850
Title:       Iter Vehems ad Necem
Description: Ett grafiskt rogue-liknande spel.
End
