Begin3
Language:    SV, 850
Title:       Ranish Partition Manager
Description: Partition Manager kan: spara och �terst�lla MBR; skapa och ta bort partitioner; visa en h�rddisks IDE-information; formatera och �ndra storlek p� FAT-16 och FAT-32 filsystem; en avancerad uppstartshanterare medf�ljer.
Keywords:    disk, partition, hanterare, ranish, fdisk, format
End
