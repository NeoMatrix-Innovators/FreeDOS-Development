Begin3
Language:    SV, 850
Title:       NGE Nibbles
Description: En klon av Nibbles, ett gammalt arkadspel.
Keywords:    nibbles
End
