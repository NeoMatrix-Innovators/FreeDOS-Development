FD-REPOv1	Build time: 1645361091	Arkivprogram	11
7zdec	17.00 beta (rev A)	uppackare f�r .7z-filer	6c57d9b1
arj	2.78a	ARJ-arkivprogrammet med �ppen k�lkod.	ed591315
bz2	1.0.8a	BZIP2-kompressionprogram	47c8c90c
cabext	1.8a	CABExtract kan extrahera filer fr�n en m�ngd olika Microsoft CAB-format.	357ee2a5
gzip	1.2.4a	GNU zip-komprimering - ett filarkvieringsverktyg, i stil med PKZIP	5e2d3f37
lpq1	2a	lpq1 �r en filkomprimerare och arkivprogram	070fc1b4
p7zip	4.65a	p7zip �r en snabb portering av 7za.exe (kommandoradsversionen av 7zip). 7-Zip �r ett filarkveringsprogram med den h�gsta kompressiongraden.	81c055e7
tar	1.12a	Ett arkivprogram f�r kassett	f90e739d
unzip	6.00a	Ett fildekomprimeringsverktyg i stil med PKUNZIP.	0a8a4d72
zip	3.0	Ett filarkivprogram i stil med PKZIP.	7efefc96
zoo	2.1a	Manipulera zoo-arkiv.	5948a9c2
