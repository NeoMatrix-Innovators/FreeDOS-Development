Begin3
Language:    SV, 850
Title:       FDTUI
Description: Text-gr�nssnitskal f�r FreeDOS
Keywords:    freedos, skal
End
