Begin3
Language:    SV, 850
Title:       FancyMines
Description: En minr�jliknande spel med snygg grafik.
Keywords:    mines
End
