Begin3
Language:    SV, 850
Title:       Blocek
Description: En grafisk textredigerare med st�d f�r unicode och bildformat
Keywords:    redigerare, unicode
End
