Begin3
Language:    SV, 850
Title:       DOSHEXED
Description: Hex-redigerare och -visare
Keywords:    hex-redigerare visare fels�kning
End
