Begin3
Language:    SV, 850
Title:       ETHTOOLS
Description: En upps�ttning diagnostikverktyg f�r ethernet-n�tverkt. Byggt med hj�lp av WatTCP-stacken. Inkluderar ETHWHAT, WWWATCH, ETHSEND, ETHDUMP, ETHWATCH, ETSHOW,
Keywords:    ethtools
End
