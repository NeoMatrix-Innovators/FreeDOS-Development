Begin3
Language:    SV, 850
Title:       LPT-drivrutin
Description: Ett verktyg f�r att styra LPT-anslutna enheter manuellt eller p� tidsbasis
Keywords:    LPT
End
