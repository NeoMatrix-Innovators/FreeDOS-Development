Begin3
Language:    SV, 850
Title:       Bolitaire
Description: En DOS-klon av Freecel 
End
