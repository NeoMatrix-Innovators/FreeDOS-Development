Begin3
Language:    SV, 850
Title:       CHKDSK
Description: Kontrollera disken efter fel.
Keywords:    kontrollera diskfel
End
