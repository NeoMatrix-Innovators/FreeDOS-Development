Begin3
Language:    SV, 850
Title:       Freedoom
Description: SMMU �r en Doom-k�llkodsportering baserad p� MBF och Boom. Denna versoin �r paketerad med Freedoom f�r en komplett spelupplevelse.
Keywords:    doom, boom, Freedoom
End
