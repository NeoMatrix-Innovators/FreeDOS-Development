Begin3
Language:    SV, 850
Title:       WDE
Description: Wde �r en diskredigerare.
Keywords:    Wde, disk, redigerare
End
