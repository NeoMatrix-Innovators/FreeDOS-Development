Begin3
Language:    SV, 850
Title:       Defrag
Description: Defragmenteringsverktyg.
Keywords:    defragmenterare
End
