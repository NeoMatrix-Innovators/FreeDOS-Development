FD-REPOv1	Build time: 1645361091	Spel	28
bolitare	0.62b	En DOS-klon av Freecel	224feeb6
boom	2.02a	En GPL-portering av Doom-k�llkoden. Paketerad med FreeDoom f�r att f� en komplett spelupplevelse.	5dbc91d6
dosdef	1.00a	DOS Defender �r ett x86 Real Mode-spel f�r DOS f�r Ludum Dare #31 (December, 2014). Eftersom endas ett f�tal DOS-maskiner fortfarande existerar �r m�lplattformen egentligen DOSBox, men det b�r fungera i viss utstr�ckning p� vilket DOS-system som helst. Spelet kan spelas med musen men �r avsett att spelas med en joystick/spelkontroll.	d61ee06b
eliza	1.01a	En av de tidigaste datorbaserade AI-tjattrobotarna	f9850151
empong	0.91a	Emeritus Pong �r en klong av det gamla h�rliga spelet Pong.	52985e35
ev4de	1.2a	EV4DE (uttalas 'ev�jd') �r ett spel om att flyga ett skepp genom rymden och undvika asteroider. Spela i tre olika spelll�gen, l�s upp ytterligare skepp och f� h�gsta po�ng! EV4DE kan spelas med ett tangentbord, men jag rekommenderar starkt att anv�nda en joystick eller spelkontroll.	3b6610b9
ewsnake	0.5a	En klon av det klassiska ormspelet (ocks� k�nt som nibbles).	23a4dbe0
flpybird	1.0a	Floppy Bird �r en klon av det �k�nda Flappy Bird skriven i 16 -bitars (x86) assembler. Med andra or fungerar det p� RENT KISEL och kr�ver inte ett underliggande operativsystem, det �r ett operativsystem i sig.	ad292fd8
fmines	1.00a	En minr�jliknande spel med snygg grafik.	6a56b580
freedoom	3.30b	SMMU �r en Doom-k�llkodsportering baserad p� MBF och Boom. Denna versoin �r paketerad med Freedoom f�r en komplett spelupplevelse.	85fb87e3
gnuchess	4.0 patch 60 (rev A)	GNU Chess �r ett gemensamt schackprogram. Bidragsgivare donerar sin tid och anstr�nging f�r att g�ra det till ett starkare, b�ttre och elegantare program.	46f36a97
hangman	1.05b	Flerspr�kig h�nga gubben	b173eadd
ivan	0.50a	Ett grafiskt rogue-liknande spel.	4f6b5e97
kraptor	Apr_2004 (rev A)	Kraptor �r ett Raptor-liknande spel med �ppen k�llkod, komplett med flera banor.	b36aaf4b
liquiwar	5.6.3a	Ett unikt krigsspel f�r flera spelare.	5401d9b0
mirmagic	2.0.2a	Ett spel i arkadstil likt Deflektor (C 64) eller Mindbender (Amiga)	94e0c875
mistral	1.0	Ett retro-RPG med spiontema och rundor f�r din klassiska maskin.	beb32643
nethack	3.4.3a	Ett spel f�r en spelare som utforskar en grotta.	d104b799
nge_nibb	0.1.0a	En klon av Nibbles, ett gammalt arkadspel.	a2200bf9
noudar	1.2	F�rsta-persons grottkravlare, anv�nder programvarurendering och fixpunktsmatte	f71896d2
qtetris	1.4.1a	En klon av spelet TETRIS, och p� samma g�ng en hyllning till bandet Queen.	b017ab63
senet	1.0a	Ett mycket gamalt spel som daterar tillbaka till forntida Egypten	3c5bee15
smiley	2021-11-10 alpha	Ett enkelt spel i pong-stil (VGA, 386+)	a8feccfa
sudoku86	1.0.3a	Ett 16-bitars Sudoku-spel f�r DOS och 8086/8088 CPU:er	9e0d8f33
vertigo	0.26a	Flygsimulator som fokuserar p� realism i flygmodellen.	10627770
vitetris	0.55a	En terminal-baserad Tetris-klon.	c303363a
wing	0.7a	Ett galaga-liknanan rymdskjutspel.	31da5be0
zmiy	0.85.2a	Ett ormspel (likt Nibbles) f�r DOS och 8086	1ad03ce9
