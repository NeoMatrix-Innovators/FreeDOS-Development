Begin3
Language:    SV, 850
Title:       ANSiMat
Description: ANSiMat �r en grafisk visare f�r ANSI-filer. Den kan ocks� anv�ndas f�r att konvertera ANSI-filer till vanliga grafikfiler (BMP/PCX/PPM/TGA/TIF) eller FLiC-animationer (FLC.
Keywords:    ansi, visare
End
