Begin3
Language:    SV, 850
Title:       NTOOL
Description: NTOOL �r ytterligare en inkarnation av det ber�mda programmet NETCAT, baserad p� WatTCP-stacken.
Keywords:    ntool,netcat
End
