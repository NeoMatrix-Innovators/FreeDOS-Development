Begin3
Language:    SV, 850
Title:       FoxCalc
Description: En snygg kalkylator. En har ett textgr�nssnit och musst�d.
Keywords:    kalkyl, FoxCalc, kalkylator, FreeDOS, Fox
End
