Begin3
Language:    SV, 850
Title:       MPlayer
Description: MPlayer �r en videospelare porterad fr�n Linux.
Keywords:    multimedia,grafik,spelare
End
