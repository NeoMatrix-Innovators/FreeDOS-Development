Begin3
Language:    SV, 850
Title:       OSPlus Text Editor
Description: En v�nlig textredigerare f�r DOS
Summary:     OSPlus Textredigerare: En v�nlig textredigrerare f�r DOS. Inkluderar Real och Protected mode-versioner (DJGPP).
Keywords:    text, redigerare, dos, rtf, txt, wri
End
