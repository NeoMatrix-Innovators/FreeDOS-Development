Begin3
Language:    SV, 850
Title:       zmiy
Description: Ett ormspel (likt Nibbles) f�r DOS och 8086
Keywords:    nibbles, snake
End
