Begin3
Language:    SV, 850
Title:       elvis
Description: En klon av vi/ex, UNIX standardredigerare. Har st�d f�r n�stan alla vi-/ex-kommandon
Keywords:    vi, redigerare
End
