Begin3
Language:    SV, 850
Title:       Dungeons of Noudar 3D
Description: F�rsta-persons grottkravlare, anv�nder programvarurendering och fixpunktsmatte
Summary:     En f�rstapersons 2.5D grottutforskare f�r Protected Mode, skrivet i C++14 (ungef�r) som ett k�rleksbrev till 90-talets RPG:er. Ljudalternativ inkluderar Adlib, PC-h�gtalare och OPL2LPT.
Keywords:    spel, rpg
End
