Begin3
Language:    SV, 850
Title:       FindDisk
Description: Litet verktyg f�r att hitta en diskett efter etikett
Keywords:    freedos, disk
End
