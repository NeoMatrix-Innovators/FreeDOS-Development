Begin3
Language:    SV, 850
Title:       TDE (Thomson-Davis Editor)
Description: TDE �r en enkel bin�r-/textfilsredigerare f�r flera filer/f�nster skriven f�r IBM PC och kompatibler som k�r DOS, Win32 (konsol)
Keywords:    redigera, redigerare, text
End
