Begin3
Language:    SV, 850
Title:       Bootfix
Description: Bootfix �r ett test- och fixverktyg f�r startsektorer.
Keywords:    Bootfix, uppstart, sektor, mbr, disk
End
