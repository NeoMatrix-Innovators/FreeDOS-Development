Begin3
Language:    SV, 850
Title:       Dialog
Description: Visa dialogrutor i skalskript
Keywords:    dialog, curses
End
