Begin3
Language:    SV, 850
Title:       Flashrom
Description: Generellt eeprom-fastprogramvara och s�kerhets-/uppdateringsverktyg f�r BIOS
Keywords:    flashrom flash bios fastprogramvara uefi efi
End
