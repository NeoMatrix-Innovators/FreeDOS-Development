Begin3
Language:    SV, 850
Title:       EW Snake
Description: En klon av det klassiska ormspelet (ocks� k�nt som nibbles).
Keywords:    snake, nibble
End
