Begin3
Language:    SV, 850
Title:       utf8tocp
Description: Konverterar UTF-8 textfiler till andra kodsidor och tillbaka
Keywords:    kodsida,konverterare
End
