FD-REPOv1	Build time: 1645361091	Applikationer	7
dn2	2.14 beta (rev A)	DOS Navigator 2 �ppen k�llkod�r en filhanterare baserad p� DOS Navigator (c) 1991-99 av RIT Research Labs.	38c2aa4f
doszip	2.55b	En liten LFN-medveten filhanterare med inbyggd zip-uppackare. Den �r byggd med JWasm och OpenWatcom. Inkluderar fullst�ndig k�llkod f�r DOS och Windows	1621b0c1
fdimples	0.11.5	FreeDOS installationsprogram - min programvara f�r paketlistredigering	592db6ed
fdshell	0.10beta (rev B)	DOSSHELL grafiskt anv�ndargr�nssnit implementerat f�r FreeDOS	972b868b
fdtui	0.8	Text-gr�nssnitskal f�r FreeDOS	d0196837
imgedit	2022-02-10 alpha	Enkle bildredigerare	4cbc3e5f
pgme	2022-02-08	En fullt konfigurerbar programstartare med flera menyer f�r DOS. Det inkluderar ocks� Font Designer och flera andra verktyg. (Kr�ver mus)	dd323bb0
