Begin3
Language:    SV, 850
Title:       CABExtract
Description: CABExtract kan extrahera filer fr�n en m�ngd olika Microsoft CAB-format.
Keywords:    cab, komprimerat, arkiv
End
