Begin3
Language:    SV, 850
Title:       TETRIS Queen
Description: En klon av spelet TETRIS, och p� samma g�ng en hyllning till bandet Queen.
Keywords:    tetris
End
