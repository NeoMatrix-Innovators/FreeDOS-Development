Begin3
Language:    SV, 850
Title:       shext
Description: Share Extender
Keywords:    delning ut�kning
End
