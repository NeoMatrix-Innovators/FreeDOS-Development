Begin3
Language:    SV, 850
Title:       FreePascal
Description: En 32-/64-bitars Pascal-kompilator som kan kompilera sig sj�lv med st�d f�r Turbo- och Delphi-dialekter. (Delar kr�ver LFN-st�d)
Keywords:    pascal, programmering, kompilator
End
