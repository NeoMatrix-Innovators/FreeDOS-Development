Begin3
Language:    SV, 850
Title:       FoxType
Description: Avancerad textfilsvisare med st�d f�r UTF-8
Keywords:    text, visare, UTF-8, UTF8, Unicode, DOS
End
