Begin3
Language:    SV, 850
Title:       rawrite
Description: Skriver diskfiler till r�a disketter
Keywords:    diskett, skriv, rawrite
End
