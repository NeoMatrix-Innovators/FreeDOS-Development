Begin3
Language:    SV, 850
Title:       EDLIN
Description: Programmet edlin �r FreeDOS standard rad-redigerare. (UPX-komprimerad)
Keywords:    redigera, redigerare, radredigerare
End
