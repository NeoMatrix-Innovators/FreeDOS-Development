FD-REPOv1	Build time: 1645361091	FreeDOS Bas	57
ambhelp	0.1d	FreeDOS-hj�lpfiler i AMB -ormat	d9c00480
append	5.0-0.6a	APPEND l�ter program �ppna datafiler i angivna kataloger som om de befanns sig i den aktuella katalogen.	882e3330
assign	1.4a	Tilldela en enhetsbokstav till en annan enhet	ba3ce6a3
attrib	2.1a	Visa och s�tt filattribut	ae4c81af
chkdsk	beta 0.9.2 (rev A)	Kontrollera disken efter fel.	06ae0e52
choice	4.4a	Presentera ett alternativ f�r anv�ndaren och v�nta p� en tangent (anv�nder kitte ist�llet f�r cats)	dccfb443
comp	1.04a	J�mf�r filer och visa deras skillnader	11355af9
cpidos	3.0a	Paket DISPLAY-typ, UPX-komprimerade CPI-filer f�r diverse DOS-kodsidor.	403e3184
ctmouse	2.1b4	FreeDOS musdrivrutin	835c58f7
debug	1.28pre1	Ett verktyg f�r programtestning och redigering	53f0f08d
defrag	1.3.2a	Defragmenteringsverktyg.	326adc6a
deltree	1.02g.mrlg (rev A)	Ta bort filer och kataloger med all inkluderade filer och underkataloger!	740f2021
devload	3.25a	Inl�sningprogram f�r drivrutiner p� kommandoraden, har st�d f�r UMB:er	6380b1c1
diskcomp	06jun2003 (rev A)	Diskj�mf�reelseverktyg	37609f47
diskcopy	beta 0.95 (rev A)	Kopiera en disk eller avbildningsfil till en annan	abba59db
display	0.13d	FreeDOS drivrutin f�r kodsideshantering (sk�rm eller skrivare)	3775e005
edit	0.9b	FreeDOS f�rb�ttrad klon av MS-DOS Edit	88e24f30
edlin	2.19	Programmet edlin �r FreeDOS standard rad-redigerare. (UPX-komprimerad)	bdcba7a1
exe2bin	1.5a	Konvertera en exe-fil till bin-format	85755cd8
fc	3.03a	Filj�mf�relseverktyg	2c92bcc7
fdapm	2009sep11 (rev A)	APM/ACPI styrning/info, str�mspar TSR/styrning, cachet�mning, omstart... {en ers�ttare f�r MS-DOS POWER}	ea7b5973
fdhelper	1.3.5	Kommandofiler f�r att utf�ra diverse uppgifter i FreeDOS	4443ed62
fdisk	1.3.4a	Verktyg f�r fixa diskar - skapa partitioner.	fb8da4c6
fdxms286	0.03.Temperaments (rev A)	Ers�ttnings-drivrutin f�r XMS f�r '286-system eller b�ttre.	66b09d32
fdxms	0.94.Bananas (rev A)	Ers�ttnings-drivrutin f�r XMS f�r '386-system eller b�ttre	aecab5d7
find	3.0b LFN (rev A)	Visa alla rader i en eller flera filer som inneh�ller en given str�ng. Omv�nda och skiftl�gesok�nsliga s�kningar ocks� m�jliga.	f5f878b4
format	0.91x	Diskformateringsprogram -- skapar FAT-filsystem och l�gniv�formaterar disketter	5deb28c4
freecom	0.85a	FreeDOS kommandoskal	f826a7c3
graphics	2008-07-14a	Till�t Prtscr att skriva ut grafiksk�rmar. (CGA/EGA/VGA/MCGA p� Postskript, ESC/P Epson 8/24-n�lars- och HP PCL-skrivare)	acd9ab1f
himemx	3.36	HimemX �r en XMS-minneshanterar baserade p� FreeDOS Himem.	931e9d67
htmlhelp	1.0.8b	HTML-visare och inneh�ll f�r FreeDOS-hj�lp	7c4da3bc
jemm	5.79d	Jemm386 �r en expanderad minneshanterare f�r DOS	5e6c77c9
kernel	2043	FreeDOS-k�rnan	128a5a03
keyb_lay	3.1a	Tangentbordslayouter f�r KEYB	f2863a2a
keyb	2.01a	Tangentbordsdrivrutin (BIOS-niv�) f�r internationellt st�d	f9cb5546
label	1.5	S�tter eller �ndrar diskens volymetikett	360f8d35
lbacache	2009feb06	Diskcache, cachar l�sningar f�r upp till 8 CHS/LBA-h�rddiskar och disketter. XMS, 386 eller b�ttre - lbacache f�ljer med tickle!	623b2399
mem	1.11a	Visar m�ngden anv�nt och fritt minne i ditt system	e0a37ac5
mirror	0.2a	Spelar in information om disken f�r eventuellt data�terst�llning.	53ebe07f
mkeyb	0.46	V�ldigt liten tangentbordsdrivrutin, 500-700 byte resident	0e64ed5f
mode	2015-11-25a	S�tt l�get f�r dina enheter:	a1378dbb
more	4.3a	Visar inneh�llet i en textfil en sida �t g�ngen	23c9b00d
move	3.3b	Flyttar filer h�rifr�n till dit	2adecd5f
nansi	4.0d (2007may26) (rev A)	En ANSI-drivrutin f�r DOS	8359ea54
nlsfunc	0.4a	NLSFUNC l�gger till NLS-funktionalitet (Nationellt spr�kst�d)	d0c3d660
print	1.02.ea (rev A)	Skriv ut filer i bakgrunden medan du g�r andra saker.	4304f677
recover	0.1 (BETA) (rev A)	�terst�ller diskar eller f�rlorad filer.	4690837c
replace	1.2a	Ers�tter filer i destinationskatalogen med filer fr�n k�llkatalogen som har samma namn.	fad75d24
samcfg	20110719a	En upps�ttning av exempelfiler f�r att skapa C:CONFIG.SYS och C:AUTOEXEC.BAT	ce19ae9e
share	08/2006a	Installerar fildelning och l�sningsm�jligheter p� din h�rddisk - endast f�r FreeDOS-k�rnan	a548904b
shsucdx	3.08a	En fri CDROM-extender f�r DOS	18d2f4f6
sort	1.5.1a	Sortera inneh�llet i en textfil, sortera valfritt enligt NLS-tabell	143218e9
swsubst	3.2a	SUBST och JOIN	5a2ead3b
tree	3.7.2a	Visar katalogstrukturen grafiskt f�r en enhet eller s�kv�g.	73317948
undelete	2008a	Undelete l�ter dig �terst�lla borttagna (men �terst�llbara) filer fr�n FAT16/FAT32-filsystem.	0230392b
unformat	0.8a	Unformat kan �terst�lla en disk som du formaterat av misstag.	4112be1d
xcopy	1.4a	Kopierar filer och katalogstr�d.	bf4ae60a
