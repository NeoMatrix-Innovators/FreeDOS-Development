FD-REPOv1	Build time: 1645361091	N�tverk	31
arachne	1.99	en webbl�sare f�r DOS (8086- & i386-versioner)	fa0d73e3
crynwr	2006-09-02c	En samling av fria paketdrivrutiner fr�n f�retaget Crynwr	e375b46d
curl	7.77.0	Curl �r ett kommandoradsverktyg f�r att �verf�ra data angiven med URL-syntax.	e0b7c5a1
dillo	3.0p9a (rev B)	En grafisk webbl�sare k�nd f�r sin hastighet och lilla minnesavtryck.	df849702
dwol	1.0a	Ett litet verktyg som ber�knar och skickar wake-on-lan-paket	322dfd21
e1000pkt	February 1, 2007 (rev A)	Paketdrivrutin f�r Intel(R) PRO/1000-kort, t.ex. 82544-, 82540-, 82545-, 82541- och 82547-baserade Ethernet kontrollerkort.	806489aa
e100pkt	0.2a	Paketdrivrutin f�r DOS	141af3c6
etherdfs	0.8.2a	Ethernet DOS-filsystem (mappare en fj�rrenhet �ver r� Ethernet)	2c7e5118
ethtools	8feb2010 (rev A)	En upps�ttning diagnostikverktyg f�r ethernet-n�tverkt. Byggt med hj�lp av WatTCP-stacken. Inkluderar ETHWHAT, WWWATCH, ETHSEND, ETHDUMP, ETHWATCH, ETSHOW,	fde3a0c2
fdnet	2022-01-11	Paket f�r grundl�ggande n�tverksst�d f�r FreeDOS. (baserat p� Rugxulos MetaDOS)	6650e592
gopherus	1.2a	En fri, (16-bitars) konsolll�gesklient f�r gopher f�r flera plattformar	bbe5c905
htget	1.06a	HTGET �r en filh�mtare som h�mtar filer fr�n HTTP-servrar.	2155309a
links	2.25	Links �r en Lynx-liknande text och grafisk WWW-l�sare.	581cb740
lsppp	1.0	En liten DOS PPP-paketdrivrutin	20c6a2b7
lynx	2.9.0-dev.10r2	Lynx text och grafik WWW-l�sare (DJGPP-portering)	958baffb
m2wat	0.1a	Verktyg f�r att �verf�ra inst�llningar fr�n MTCP.CFG till WATTCP.CFG.	d6568304
mskermit	3.16a	Kommunikationssvit fr�n Columbia universitetet.	0b7491f9
mtcp	2020-03-07	En UPX:ad samling TCP/IP-verktyg f�r 16-bitars DOS: DHCP, IRC, FTP, Telnet, Netcat, HTGet, Ping, SNTP	6c876606
newsnuz	0.98a	Usenet-l�sare (NNTP) baserad p� WatTCP	21ce4a27
ntool	1.5a	NTOOL �r ytterligare en inkarnation av det ber�mda programmet NETCAT, baserad p� WatTCP-stacken.	e6f4a6db
picosntp	0.9.1a	SNTP-klient f�r DOS, baserad p� picoTCP	fd13e8eb
picotcp	20151119a	picoTCP-n�tverksstack (bibliotek och konfigurationsverktyg)	63458220
ping	2.2a	Verktyget ping f�r internetdiagnostik. Denna version extraherades fr�n Watt-32 v2.2-sviten.	35b92e05
rsync	2.2.5a	rsync �r en verktygsprogramvara som synkroniserar filer och kataloger fr�n en plats til en annan medan det minimerar data�verf�ring genom deltakodning n�r s� �r l�mpligt. Denna rsync-portering �r n�dv�ndigtvis en delm�ngd av den fulla rsync, delvis p� grund av minnebegr�nsningar och delvis p� grund av egenheter hos DOS. Huvudskillnaderna �r: Endast f�r klient; inget st�d f�r rsh eller ssh; filnamn p� servern m�ste vara i DOS-format; fildata komprimeras inte.	2ae9d57f
ssh2dos	0.2.1a	SSH-klient f�r SSH-protokoll version 2.0. Inneh�ller ocks� SCP, SFTP och telnet i b�de 8086- och 386-versioner.	8b129854
sshdos	0.95a	SSH-klient f�r DOS. Inneh�ller ocks� SSH, SCP och SFTP i b�de 8086- och 386-versioner.	84b2ae5a
terminal	3.2a	En liten vt100/ansi-terminale f�r varje pc	85f77c4a
vmsmount	0.5c	En DOS-omdirigerare f�r montering av VMware:s delade mappar	9cf80608
vncview	3.3.7a	VNC-visare f�r 8086+, baserad p� Xvncviewer	dde4b5b9
wattcp	2016-05-19a	WATTCP	fa7b5ade
wget	1.11.2a	Icke-interaktiv n�tverksh�mtare.	1598769b
