Begin3
Language:    SV, 850
Title:       ETHERDFS
Description: Ethernet DOS-filsystem (mappare en fj�rrenhet �ver r� Ethernet)
Summary:     EtherDFS �r en 'installerbart filsystem'-TSR f�r DOS. Det mappar en enhet fr�n en fj�rrdator (typiskt Linux-baserad) till en lokal enhetsbokstav, som anv�nder r�da ethernetpaket f�r att kommunicera. Under m�nga �r anv�nde jag LapLink f�r att �verf�ra filer mellan alla mina retrodatorer. Ja, det fungerar men det �r ocks� irriterande l�ngsamt och kr�ver konstant uppm�rksamhet. On dag t�nkte jag: 'Vore det inte fantastiskt om alla mina DOS PC kunde dela en gemensam n�tverksenhet, liknande hur NFS fungerar i *nix-v�rlden?'. Den dagen f�ddes EtherDFS. Jag har helt klart inte uppfunnit n�got - konceptet har funnit n�stan lika l�nge som den f�rsta IBM PC:n, och flera kommersiella produkter har adresserat detta behovet tidigare. Men jag k�nner inte till n�gon fri l�sning med �ppen k�llkod. Dessutom kr�ver alla kommersiella l�sningar jag k�nner till att du f�rst s�tter upp en ganska komplicerad n�tverksmilj�, medan EtherDFS inte kr�ver n�got mer �n en paketdrivrutin.
Keywords:    etherdfs
End
