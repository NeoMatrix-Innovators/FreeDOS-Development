FD-REPOv1	Build time: 1645361091	Utveckling	6
bcc	0.16.10a	Bruce's C compiler �r en enkel C-kompilator som producerar 8086-assembler f�r minnesmodellerna tiny/small.	7bed01aa
fpc	3.2.2	En 32-/64-bitars Pascal-kompilator som kan kompilera sig sj�lv med st�d f�r Turbo- och Delphi-dialekter. (Delar kr�ver LFN-st�d)	1bb88014
kittenc	2021-08-01	catgets/kittengets-kompatibel resurskompilator	c4fbf05d
nasm	2.15.05a	Netwide Assembler (UPX-komprimerad version)	b33948e8
upx	3.96a	UPX �r ett fritt, portabelt, ut�kningsbart, h�gpresterande kompressionprogram f�r k�rbara filer f�r m�nga olika format.	be14f7f2
watcomc	1.9	Open Watcom C-/C++-kompilator	9c22f267
