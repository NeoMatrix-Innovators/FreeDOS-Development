Begin3
Language:    SV, 850
Title:       DOS/32A
Description: DOS/32A �r en DOS extender.
Keywords:    7-zip, 7z, 7za, arkivprogram
End
