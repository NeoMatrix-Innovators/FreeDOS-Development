Begin3
Language:    SV, 850
Title:       PRINT
Description: Skriv ut filer i bakgrunden medan du g�r andra saker.
Keywords:    skriv ut, spooler, lpr
End
