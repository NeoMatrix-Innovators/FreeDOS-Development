Begin3
Language:    SV, 850
Title:       TAR (GNU TAR)
Description: Ett arkivprogram f�r kassett
Keywords:    arkivprogram, kassett
End
