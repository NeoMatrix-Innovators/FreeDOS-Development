Begin3
Language:    SV, 850
Title:       Vi IMproved (vim)
Description: F�rb�ttrad version av textredigeraren vi.
Summary:     VIM �r en f�rb�ttrad version av redigeraren vi, en av standardtextredigerarna p� UNIX-system. Dessa �r k�rtidsfiler f�r VIM. [GPL-kompatibel, men om du tycker att det �r anv�ndbart ber dig g�ra en donation f�r att hj�lpa barn i Uganda via ICCF. Den fullst�ndiga licenstexten kan hittas i README.txt.] Endast 32-bitars dos (sedan 7.1).
Keywords:    redigerare, vi, vim
End
