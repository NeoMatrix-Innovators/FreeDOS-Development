Begin3
Language:    SV, 850
Title:       KEYB layouter
Description: Tangentbordslayouter f�r KEYB
Keywords:    keyb,layouter
End
