Begin3
Language:    SV, 850
Title:       nro
Description: En textbehandlare i stil med nroff i UNIX
Keywords:    nroff, roff, nro, micro-c
End
