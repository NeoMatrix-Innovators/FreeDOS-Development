Begin3
Language:    SV, 850
Title:       SSHDOS
Description: SSH-klient f�r DOS. Inneh�ller ocks� SSH, SCP och SFTP i b�de 8086- och 386-versioner.
Keywords:    ssh protokoll n�tverk kommunikation fj�rr�tkomst
End
