Begin3
Language:    SV, 850
Title:       Localize
Description: �vers�tter texter
Keywords:    freedos lokalisera kommandofil
End
