Begin3
Language:    SV, 850
Title:       The Mistral Report: Invisible Affairs
Description: Ett retro-RPG med spiontema och rundor f�r din klassiska maskin.
Summary:     The Mistral Report: Invisible Affairs �r ett retro-RPG med spiontema baerat p� rundor f�r din klassiska maskin. Kr�ver 386SX eller b�ttre. Ljudalternativ inkluderar Adlib, PC-h�gtalare och OPL2LPT.
Keywords:    spel, rpg
End
