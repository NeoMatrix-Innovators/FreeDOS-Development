Begin3
Language:    SV, 850
Title:       Boom
Description: En GPL-portering av Doom-k�llkoden. Paketerad med FreeDoom f�r att f� en komplett spelupplevelse.
Keywords:    doom,boom,freedoom
End
