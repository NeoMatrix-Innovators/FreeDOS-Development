Begin3
Language:    SV, 850
Title:       Syslinux
Description: Syslinux samling av uppstartsprogram
Keywords:    eltorito syslinux memdisk isolinux modulkedja
End
