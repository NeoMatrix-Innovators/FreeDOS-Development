Begin3
Language:    SV, 850
Title:       DOSFSCK
Description: Kontrollerar PC/MS-DOS filsystem och f�rs�ker valfritt reparera dem
Keywords:    scandisk,chkdsk
End
