Begin3
Language:    SV, 850
Title:       Wget
Description: Icke-interaktiv n�tverksh�mtare.
Keywords:    freedos, wget
End
