Begin3
Language:    SV, 850
Title:       PG (PaGer)
Description: Visar inneh�llet i en textfil en sida �t g�ngen
Keywords:    sida, text, visa text
End
