Begin3
Language:    SV, 850
Title:       SetLock
Description: St�ller in Caps-, Num- och Scroll-lock-tangenterna fr�n programvara
Keywords:    l�s, caps, num, scroll, s�tt
End
