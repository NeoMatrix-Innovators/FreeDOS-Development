Begin3
Language:    SV, 850
Title:       XGREP
Description: Snabb UNIX-liknande `grep'-klon med st�d f�r regulj�ra uttryck
Keywords:    freedos, filer, hitta, grep, s�k, text, unix-like
End
