Begin3
Language:    SV, 850
Title:       Open Watcom C-kompilator
Description: Open Watcom C-/C++-kompilator
Keywords:    watcom, c, kompilator
End
