Begin3
Language:    SV, 850
Title:       Callver
Description: S�tter DOS-versionen under ett programs k�rning.
Keywords:    Dos FreeDOS setver dosver callver version
End
