Begin3
Language:    SV, 850
Title:       DELTREE
Description: Ta bort filer och kataloger med all inkluderade filer och underkataloger!
Keywords:    freedos, ta bort, tr�d
End
