Begin3
Language:    SV, 850
Title:       LSppp
Description: En liten DOS PPP-paketdrivrutin
Keywords:    paket
End
