Begin3
Language:    SV, 850
Title:       CDP
Description: Audio CD-spelare f�r DOS kommandorad
Keywords:    cdp, ljud, cd-rom
End
