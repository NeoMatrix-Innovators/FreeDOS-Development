Begin3
Language:    SV, 850
Title:       picoSNTP
Description: SNTP-klient f�r DOS, baserad p� picoTCP
Keywords:    NTP, SNTP
End
