Begin3
Language:    SV, 850
Title:       AMB Reader
Description: l�sare f�r Ancient Machine Book-formatet
Summary:     AMB �r en l�sare f�r AMB-filer, som st�r f�r Ancient Machine Book. Det �r ett extremt l�ttviktigt filformat menat f�r att spara alla typer av hypertext-dokument som bekv�mt kan l�sas p� �ven de mest forntida datorerna: tekniska manualer, b�cker, osv. T�nk p� det som en retro-variant av en *.CHM-hj�lpfil.
Keywords:    text, dokument, l�sare
End
