Begin3
Language:    SV, 850
Title:       freemacs
Description: En emacs-liknande redigarare f�r DOS (likt GNU Emacs)
Keywords:    redigera, redigerare, unicode
End
