Begin3
Language:    SV, 850
Title:       7zdec
Description: uppackare f�r .7z-filer
Summary:     listen, frist�ende dekomprimerare f�r 7-Zip-arkiv (med ANSI C-k�llkod)
Keywords:    7z, 7zdec, 7zdecode, arkiv
End
