Begin3
Language:    SV, 850
Title:       GNU Chess
Description: GNU Chess �r ett gemensamt schackprogram. Bidragsgivare donerar sin tid och anstr�nging f�r att g�ra det till ett starkare, b�ttre och elegantare program.
Keywords:    chess,gnuchess
End
