FD-REPOv1	Build time: 1645361091	Verktyg	56
aefdisk	1.0a	Kommandoradsdrivet diskpartitioneringsverktyg f�r DOS (portat f�r Open Watcom)	fe87ee00
ambread	20201223	l�sare f�r Ancient Machine Book-formatet	3845698b
ansimat	0.93a	ANSiMat �r en grafisk visare f�r ANSI-filer. Den kan ocks� anv�ndas f�r att konvertera ANSI-filer till vanliga grafikfiler (BMP/PCX/PPM/TGA/TIF) eller FLiC-animationer (FLC.	0fd59a47
b64	0.06R (rev A)	Verktyg som implementerat Content-Transfer-Encoding-standarden Base64 beskriven i RFC1113.	f940dfeb
bmp2png	1.62a	Kommandoradsverktyg som konverterar BMP-bilder till PNG (och omv�nt)	0f396f96
bootfix	1.4a	Bootfix �r ett test- och fixverktyg f�r startsektorer.	d409f0e6
bsum	1.1a	ber�knar BSD-kontrollsummor f�r filer	2c81e33a
callver	2007-08-19a	S�tter DOS-versionen under ett programs k�rning.	b1fd312f
cdrom2ui	2003-11-16a	Ett litet verktyg f�r att mata ut, st�nga sp�ret, l�sa, l�sa upp eller �terst�lla en CD-ROM efter enhetsbokstav.	0ca5a9dd
cpied	1.3d	En GUI-driven CPI-typsnittsredigerare	dce8e6a1
cwsdpmi	7a	32-bitars DPI DOS extender designad f�r DJGPP.	68000114
dialog	1.1-20080819a	Visa dialogrutor i skalskript	5c966da5
dog	0.8.3c	Ett alternativs command.com-skal, i stil med FreeCOM, men annorlunda.	9b0fc76a
dos32a	9.1.2a	DOS/32A �r en DOS extender.	1f6e8894
dosfsck	2.11d	Kontrollerar PC/MS-DOS filsystem och f�rs�ker valfritt reparera dem	597867a7
dosutil	2012a	En samling sm� verktyg f�r kommandofiler	2d651e83
edict	0.10 (BETA) (rev A)	Enhanced Disk Image Creation Tool - ett verktyg f�r att utan problem skapa diskavbildningar f�r disketter	0c2eebaf
fdnpkg	0.99.7a	N�tverksbaserad pakethanterare	852ca0c0
finddisk	2005-03-23a	Litet verktyg f�r att hitta en diskett efter etikett	ba1f7c50
flashrom	0.9.4(-revision 1495) (rev A)	Generellt eeprom-fastprogramvara och s�kerhets-/uppdateringsverktyg f�r BIOS	eecd8007
foxcalc	0.92a	En snygg kalkylator. En har ett textgr�nssnit och musst�d.	847cedc6
foxtype	0.16a	Avancerad textfilsvisare med st�d f�r UTF-8	463a0d36
gnuchcp	1.0b	LOADFONT (GNUCHCP) �ndrar EGA-/VGA-bitmappstypsnitt p� sk�rmen i textl�ge.	f2bfcc3a
gnufonts	1.0a	LOADFONT (GNUCHCP) r�a EGA-/VGA-bitmappstypsnitt f�r textl�gen.	7552f3fd
hexcomp	1.0.4a	J�mf�r bin�rfiler grafiskt	703659ad
listpci	1.02	Visar data om PCI-enheter	5cccd490
listvesa	1.01	Verktyg f�r att rapportera vilka VESA-grafikl�gen som st�ds	77f6a43e
localcfg	0.90a	Konfigurationsverktyg f�r lokalinst�llningar	18191130
localize	1.00a	�vers�tter texter	9e837051
memteste	2003a	MEMTESTE �r ett program f�r att testa DRAM (huvudminnet) f�r PC-kompatibla datorer byggda p� Intel 386 eller senare.	45a0cce1
ospimg	1.4a	Verktyg f�r att l�sa och skriva disketavbildningar	e4cecfa1
part	2.37a	Partition Manager kan: spara och �terst�lla MBR; skapa och ta bort partitioner; visa en h�rddisks IDE-information; formatera och �ndra storlek p� FAT-16 och FAT-32 filsystem; en avancerad uppstartshanterare medf�ljer.	030a698e
pcisleep	12 mar 2005 (rev A)	PCISLEEP listar och s�ver pci-kort.	c23acedd
pdtree	1.02-1a	Visa mappstrukturen f�r en enhet eller s�kv�g grafiskt. Har st�d f�r l�nga filnamn om LFN-API:et �r installerat, st�d f�r meddelandet kataloger (olika spr�k) via cats, och st�d b�de f�r Windows NT/9x och DOS.	9f5b0a7c
pg	1.16a	Visar inneh�llet i en textfil en sida �t g�ngen	3fe5e511
pkgtools	2021-12-31	Allm�nna underh�llsverktyg f�r FreeDOS-paket	ea34f091
raread	1.1a	L�ger ut avbildningen f�r en diskett (som kan skrivas med RAWRITE). Anv�ndbart f�r att skapa diskavbildningar.	f274d322
rawrite	1.3a	Skriver diskfiler till r�a disketter	68f5edcd
rcal	1.0a	En kalkylator f�r stora tal med st�d f�r flytpunktstal som liknar pappersruller�knare. 8086+	3aa4c8ab
search	1.0a	Hittar filer p� din dator	788d1840
setlock	1.0a	St�ller in Caps-, Num- och Scroll-lock-tangenterna fr�n programvara	8119cad8
slowdown	3.10a	G�r en snabb dator l�ngsammare. Hastigheten �r helt konfigurerbar fr�n kommandoraden eller med hj�lp av snabbtangenter. Har flera olika s�tt eller l�gen f�r att g�ra datorn l�ngsammare.	05cc2a16
stamp	2.0a	S�tt, visa och filtrera tidsst�mpliar f�r filer	00deaaff
switchar	1.0a	Visa och s�tt DOS switchar	3586ba66
testdisk	7.1a	Testdisk kontrollerar partitioner/startsektorer p� diskar; Photorec �terst�ller m�nga typer av data	e796f84e
topspin	3a	Ett menytolkningsprogram som l�ger anv�ndare skapa integrerade milj�er d�r inga finns.	606ba79c
tp7p5fix	1.04	TSR f�r att att fixa fel 200 i Turbo Pascal-program vid k�rdtid utan att den k�rbara filen m�ste �ndras.	222b7ada
unrtf	0.21.5a	Konverterar dokument i RTF-format till andra format (html,latex,txt...)	0fc20871
utf8tocp	0.9.2a	Konverterar UTF-8 textfiler till andra kodsidor och tillbaka	281792ca
v8power	22.02.07	En upps�ttning av f�rb�ttringsverktyg f�r kommandofiler f�r DOS som kan tillhandah�lla textgr�nssnitt och andra behandlingsfunktioner (UPX:at)	50f478fc
wcd	6.0.2a	WCD f�r DOS byter till vilken katalog som helst, en klon av Norton Change Directory (NCD) med fler funktioner.	16fb7a22
wde	3.0c	Wde �r en diskredigerare.	b3285ecd
whichfat	2003-11-24a	K�rnst�d f�r FAT32 identifiering och FAT-typdetektering (12-32) per enhet	3963ec2f
wptail	0.52.10a	Skapa TUI-dialogruton och formul�r och samla in data fr�n anv�ndaren via libnewt	b1c631ab
xdel	2.06a	Ut�kad filborttagning, liknar DR-DOS	4e7cd24c
zerofill	1.05a	Fyller tomt utrymme p� en enhet med nollor.	435c4521
