Begin3
Language:    SV, 850
Title:       stamp
Description: S�tt, visa och filtrera tidsst�mpliar f�r filer
Keywords:    freedos
End
