Begin3
Language:    SV, 850
Title:       V8Power Tools
Description: En upps�ttning av f�rb�ttringsverktyg f�r kommandofiler f�r DOS som kan tillhandah�lla textgr�nssnitt och andra behandlingsfunktioner (UPX:at)
Keywords:    dos 16-bitars kommandofil vask vchoice vecho vpause vframe vmath vline vprogres
End
