Begin3
Language:    SV, 850
Title:       zoo
Description: Manipulera zoo-arkiv.
Keywords:    zoo
End
