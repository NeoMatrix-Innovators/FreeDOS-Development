Begin3
Language:    SV, 850
Title:       zip
Description: Ett filarkivprogram i stil med PKZIP.
Keywords:    freedos, zip, infozip, pkzip
End
