Begin3
Language:    SV, 850
Title:       trch
Description: �vers�tter tecken. Detta kan anv�ndas med programmet UNIX2DOS, men kan �vers�tta fler tecken. [Liknar, men �r inte samma som, tr i UNIX.] (inkluderar Cats GNU LGPL)
Keywords:    trch, unix2dos, tr
End
