Begin3
Language:    SV, 850
Title:       ImgEdit
Description: Enkle bildredigerare
Summary:     En enkel pixelredigerare mestadels f�r att skapa grafik f�r Danger Engine. Den har begr�nsat st�d f�r icke-inbyggda grafikformat s� som BMP. F�r n�rvaran kan vissa alternativ (s� som bildstorlek) endast st�llas in fr�n kommandoraden. Den inkluderar �ven den enkla visaren IMGVIEW. Kr�ver 386+, VGA och mus (UPX-komprimerad)
Keywords:    dos, spel, bilder, sprite:ar, igg, igs, bmp, utveckling
End
