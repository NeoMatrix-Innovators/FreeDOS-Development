Begin3
Language:    SV, 850
Title:       kittenc
Description: catgets/kittengets-kompatibel resurskompilator
Keywords:    dos, bibliotek, utveckling
End
