Begin3
Language:    SV, 850
Title:       ListVESA
Description: Verktyg f�r att rapportera vilka VESA-grafikl�gen som st�ds
Summary:     ListVESA �r ett verktyg f�r att rapportera vilka VESA-grafikl�sen som st�ds av systemets h�rdvara. Du kan anvnda kommandoradsflaggor f�r att anpass informationen som listas f�r varje l�se, l�gen soim har st�d f�r ett visst bitdjup, l�gen som har st�d f�r linj�r bildrutesbuffert eller generell information om grafikkortet i sig utan detaljerad sk�rml�gesdata.
Keywords:    lista, l�ge, VESA, grafik
End
