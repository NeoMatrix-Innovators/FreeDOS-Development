Begin3
Language:    SV, 850
Title:       OSPlus Disk Imager
Description: Verktyg f�r att l�sa och skriva disketavbildningar
Summary:     OSPlus diskavbildare �r ett verktyg som l�ter dig l�sa diskette och skapa avbildningar av dem p� din h�rddisk. Dessa kan sedan skrivas till en CD, zippas och e-postas eller skickas upp till internet. Diskavbildaren l�ter dig ocks� skriva dessa avbildningar tillbaka till en diskett. Du f�rvarnas h�r med att data p� disketten kommer att F�RST�RAS n�r du skriver en avbildning.
Keywords:    disk, avbildning
End
