Begin3
Language:    SV, 850
Title:       FDNet
Description: Paket f�r grundl�ggande n�tverksst�d f�r FreeDOS. (baserat p� Rugxulos MetaDOS)
Summary:     Tillhandah�ller grundl�ggande n�tverksst�d f�r FreeDOS p� h�rdvara/virtuella plattformar som st�ds. FDNet �r fr�n b�rjan baserat p� Rugxulo:s kommandofil CONNECT fr�n MetaDOS.
Keywords:    dos kommandofil n�tverk
End
