Begin3
Language:    SV, 850
Title:       Emeritus Pong
Description: Emeritus Pong �r en klong av det gamla h�rliga spelet Pong.
Keywords:    Pong, Spel
End
