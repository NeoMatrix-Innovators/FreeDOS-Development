Begin3
Language:    SV, 850
Title:       MEM
Description: Visar m�ngden anv�nt och fritt minne i ditt system
Keywords:    Memory, mem, xms, ems, umb, hma
End
