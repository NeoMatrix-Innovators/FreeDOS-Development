Begin3
Language:    SV, 850
Title:       rcal
Description: En kalkylator f�r stora tal med st�d f�r flytpunktstal som liknar pappersruller�knare. 8086+
Keywords:    kalkyl, kalkylator
End
