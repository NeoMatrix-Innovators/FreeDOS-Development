Begin3
Language:    SV, 850
Title:       Pico
Description: Enkel textredigerare i stil med Pine Composer
Keywords:    redigerare
End
