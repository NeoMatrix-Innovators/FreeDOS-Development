Begin3
Language:    SV, 850
Title:       ARJ
Description: ARJ-arkivprogrammet med �ppen k�lkod.
End
