Begin3
Language:    SV, 850
Title:       FDSHELL
Description: DOSSHELL grafiskt anv�ndargr�nssnit implementerat f�r FreeDOS
Keywords:    DOSSHELL GUI FreeDOS DOS
End
