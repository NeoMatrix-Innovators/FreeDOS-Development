Begin3
Language:    SV, 850
Title:       hexcomp
Description: J�mf�r bin�rfiler grafiskt
Keywords:    hex,j�mf�r
End
