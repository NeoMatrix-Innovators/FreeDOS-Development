Begin3
Language:    SV, 850
Title:       TP7/P5+-fix
Description: TSR f�r att att fixa fel 200 i Turbo Pascal-program vid k�rdtid utan att den k�rbara filen m�ste �ndras.
Keywords:    DOS, SPEL
End
