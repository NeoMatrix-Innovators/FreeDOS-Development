Begin3
Language:    SV, 850
Title:       UPX
Description: UPX �r ett fritt, portabelt, ut�kningsbart, h�gpresterande kompressionprogram f�r k�rbara filer f�r m�nga olika format.
Keywords:    komprimerare k�rbara filer
End
