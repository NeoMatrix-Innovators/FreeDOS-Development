Begin3
Language:    SV, 850
Title:       Whiptail
Description: Skapa TUI-dialogruton och formul�r och samla in data fr�n anv�ndaren via libnewt
Keywords:    dialog, whiptail, newt, gpm
End
