Begin3
Language:    SV, 850
Title:       pdTree
Description: Visa mappstrukturen f�r en enhet eller s�kv�g grafiskt. Har st�d f�r l�nga filnamn om LFN-API:et �r installerat, st�d f�r meddelandet kataloger (olika spr�k) via cats, och st�d b�de f�r Windows NT/9x och DOS.
Keywords:    tr�d, FreeDOS, DOS, Win32
End
