Begin3
Language:    SV, 850
Title:       UIDE
Description: En cachande drivrutin f�r allm�nt bruk f�r DOS-enheter, diskett, CD/DVD, SATA och UltraDMA-diskar
Keywords:    ahci, cache, cc, cd, cd-rom, cdrom, disk, dma, drivrutin, eide, diskett, ide, pata, rom, sata, sata, uhdd, uide, ultra
End
