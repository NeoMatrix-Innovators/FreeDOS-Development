Begin3
Language:    SV, 850
Title:       Eliza
Description: En av de tidigaste datorbaserade AI-tjattrobotarna
End
