Begin3
Language:    SV, 850
Title:       LFNDOS
Description: Tillhandah�ller Windows 95:s API f�r l�nga filnamn till DOS-program. DOS-program som kan anv�nda l�nga filnamn, till exempel DOS 7 Command.com, edit.com och alla DJGPP-program kan l�sa in och spara dem med hj�lp av LFNDOS. Designat f�r Win95-anv�ndare som anv�nder DOS-l�ge, men det fungerar �ven under �ldre DOS-versioner.
Keywords:    l�nga filnamn, lfn
End
