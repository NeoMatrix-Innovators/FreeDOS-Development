Begin3
Language:    SV, 850
Title:       cdrom2ui
Description: Ett litet verktyg f�r att mata ut, st�nga sp�ret, l�sa, l�sa upp eller �terst�lla en CD-ROM efter enhetsbokstav.
Keywords:    freedos, cd-rom
End
