Begin3
Language:    SV, 850
Title:       mbedit - Multi platform editor
Description: mbedit �r en helsk�rmstextredigerare med makrost�d, inbyggd kalkylator, historikbuffert f�r kommandon, hexredigerare och m�nga andra funktioner.
Keywords:    redigerare,hex
End
