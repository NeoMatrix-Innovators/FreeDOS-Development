Begin3
Language:    SV, 850
Title:       keyb
Description: Tangentbordsdrivrutin (BIOS-niv�) f�r internationellt st�d
Keywords:    keyb, tangentbord, drivrutin
End
