Begin3
Language:    SV, 850
Title:       DWOL
Description: Ett litet verktyg som ber�knar och skickar wake-on-lan-paket
Keywords:    dos n�tverk
End
