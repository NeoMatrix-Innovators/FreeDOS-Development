Begin3
Language:    SV, 850
Title:       bcc - Bruce's C compiler
Description: Bruce's C compiler �r en enkel C-kompilator som producerar 8086-assembler f�r minnesmodellerna tiny/small.
Keywords:    K&R,C89,C,kompilator
End
