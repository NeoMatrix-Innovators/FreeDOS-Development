Begin3
Language:    SV, 850
Title:       MEMTESTE
Description: MEMTESTE �r ett program f�r att testa DRAM (huvudminnet) f�r PC-kompatibla datorer byggda p� Intel 386 eller senare.
Keywords:    RAM test, memtest
End
