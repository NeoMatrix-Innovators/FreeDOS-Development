Begin3
Language:    SV, 850
Title:       less
Description: Less �r ett program i stil med more, men vilket l�ter dig g� bak�t i filen s� v�l som fram�t. Less m�ste heller inte l�sa hela indatafilen innan den startar, s� f�r st�rre indatafiler startar det upp snabbare �n textredigerare som vi.
Keywords:    less,more,sidvisare
End
