Begin3
Language:    SV, 850
Title:       EV4DE
Description: EV4DE (uttalas 'ev�jd') �r ett spel om att flyga ett skepp genom rymden och undvika asteroider. Spela i tre olika spelll�gen, l�s upp ytterligare skepp och f� h�gsta po�ng! EV4DE kan spelas med ett tangentbord, men jag rekommenderar starkt att anv�nda en joystick eller spelkontroll.
Keywords:    spel
End
