Begin3
Language:    SV, 850
Title:       EDICT
Description: Enhanced Disk Image Creation Tool - ett verktyg f�r att utan problem skapa diskavbildningar f�r disketter
Keywords:    dos 16-bitars
End
