Begin3
Language:    SV, 850
Title:       assign
Description: Tilldela en enhetsbokstav till en annan enhet
Keywords:    freedos, assign
End
