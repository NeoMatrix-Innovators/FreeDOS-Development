Begin3
Language:    SV, 850
Title:       VMSMOUNT
Description: En DOS-omdirigerare f�r montering av VMware:s delade mappar
Keywords:    vmware
End
