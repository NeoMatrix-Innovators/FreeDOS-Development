Begin3
Language:    SV, 850
Title:       LPQ1
Description: lpq1 �r en filkomprimerare och arkivprogram
Keywords:    arkivprogram, lpq1
End
