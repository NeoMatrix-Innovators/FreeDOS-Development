Begin3
Language:    SV, 850
Title:       Vitetris
Description: En terminal-baserad Tetris-klon.
End
