Begin3
Language:    SV, 850
Title:       raread
Description: L�ger ut avbildningen f�r en diskett (som kan skrivas med RAWRITE). Anv�ndbart f�r att skapa diskavbildningar.
Keywords:    r�, l�sning, diskett, avbildning
End
