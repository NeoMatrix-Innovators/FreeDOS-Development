Begin3
Language:    SV, 850
Title:       cpied
Description: En GUI-driven CPI-typsnittsredigerare
Keywords:    cpi,cpx,typsnitt,redigerare
End
