Begin3
Language:    SV, 850
Title:       ListPCI
Description: Visar data om PCI-enheter
Summary:     ListPCI �r ett verktyg f�r att list PCI-enheter som avs�ker PCI-bussen p� systemet det k�rs och visar data om alla PCI-enheter det hittar. Det tillhandah�ller mer utf�rlig data �n andra j�mf�rbara applikation och �r mer flexibelt vad det g�ller kommandoradsflaggor. Via detta kan du filtrera vilka enheter som rapporteras till att bara visa de fr�n ett specifikt tillverkar-ID eller en angiven klass. ListPCI kan ocks� returnera antalet matchande enheter i DOS-system variabel ERRORLKEVEL, vilket g�r det enkelt att integrera i kommandofiler.
Keywords:    enhet, lista, PCI
End
