Begin3
Language:    SV, 850
Title:       DOSLFN
Description: Tillhandah�ller LFN (L�nga FilNamn) API:et i ren DOS (utan Windows)
Keywords:    l�nga filnamn, lfn
End
