Begin3
Language:    SV, 850
Title:       Wing
Description: Ett galaga-liknanan rymdskjutspel.
Keywords:    galaga
End
