Begin3
Language:    SV, 850
Title:       uHex
Description: uHex �r en enkel och snabb hexredigerare
Keywords:    hex,redigerare,visare
End
