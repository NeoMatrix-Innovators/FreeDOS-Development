FD-REPOv1	Build time: 1645361091	Uppstartsverktyg	1
syslnx	4.05a	Syslinux samling av uppstartsprogram	6f7f7a6e
