Begin3
Language:    SV, 850
Title:       Vertigo
Description: Flygsimulator som fokuserar p� realism i flygmodellen.
End
