Begin3
Language:    SV, 850
Title:       HEAD
Description: Visar en del av en fil
Keywords:    head
End
