Begin3
Language:    SV, 850
Title:       wcd
Description: WCD f�r DOS byter till vilken katalog som helst, en klon av Norton Change Directory (NCD) med fler funktioner.
Keywords:    chdir, cd, �ndra katalog, snabb
End
