FD-REPOv1	Build time: 1645361091	Textredigerare	16
biew	6.10a	Biew �r en bin�r/hexadecimal visare/redigerare. (kr�ver i686+)	1fe6ebe6
blocek	1.62r2	En grafisk textredigerare med st�d f�r unicode och bildformat	c2dbe140
doshexed	1.2g	Hex-redigerare och -visare	4f1cd182
e3	2.7.1a	En liten textredigerarer som finns i b�de 32- och 16-bitars versioner	cda01462
elvis	2.2a	En klon av vi/ex, UNIX standardredigerare. Har st�d f�r n�stan alla vi-/ex-kommandon	295f17c0
fed	2.24c	En radbrytande textredigerare med f�rgmarkering av syntax och mer �n s�	a58e4e3b
freemacs	1.6h	En emacs-liknande redigarare f�r DOS (likt GNU Emacs)	59bf43d3
mbedit	8.64a	mbedit �r en helsk�rmstextredigerare med makrost�d, inbyggd kalkylator, historikbuffert f�r kommandon, hexredigerare och m�nga andra funktioner.	170f2c36
mined	2015.25a	Textredigerare med utf�rligt Unicode- och CJK-st�d. Beh�ndig och effktiva funktioner f�r redigering av rena textdokument, program, HTML, osv. Anv�ndarv�ndligt gr�nssnitt, musstyrning och menyer.	2b9519a5
msedit	0.11a	Mateusz Saucy Editor	8b351c1c
ospedit	2.1.1a	En v�nlig textredigerare f�r DOS	c9400b69
pico	3.96a	Enkel textredigerare i stil med Pine Composer	301fc35c
setedit	0.5.4a	En textredigerare f�r programmerare f�r DJGPP, liknar BC++ IDE och RHIDE	bb805916
tde	5.1w	TDE �r en enkel bin�r-/textfilsredigerare f�r flera filer/f�nster skriven f�r IBM PC och kompatibler som k�r DOS, Win32 (konsol)	6e7518af
uhex	1.0.4a	uHex �r en enkel och snabb hexredigerare	910e592c
vim	7.3a	F�rb�ttrad version av textredigeraren vi.	14cff902
