Begin3
Language:    SV, 850
Title:       VNC Viewer 8086
Description: VNC-visare f�r 8086+, baserad p� Xvncviewer
Keywords:    VNC, 8086
End
