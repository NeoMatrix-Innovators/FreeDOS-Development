Begin3
Language:    SV, 850
Title:       APPEND
Description: APPEND l�ter program �ppna datafiler i angivna kataloger som om de befanns sig i den aktuella katalogen.
Keywords:    freedos, append, data, filer, kataloger
End
