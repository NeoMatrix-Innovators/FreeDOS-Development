Begin3
Language:    SV, 850
Title:       topspin
Description: Ett menytolkningsprogram som l�ger anv�ndare skapa integrerade milj�er d�r inga finns.
Keywords:    meny, system, verktyg
End
