Begin3
Language:    SV, 850
Title:       HiRAM
Description: �vre minnesut�kare (UMB) f�r 80286, 80386, 80486 CPU:er
Keywords:    UMB,minne,hanterare
End
