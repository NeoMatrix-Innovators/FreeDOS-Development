Begin3
Language:    SV, 850
Title:       picoTCP
Description: picoTCP-n�tverksstack (bibliotek och konfigurationsverktyg)
End
