Begin3
Language:    SV, 850
Title:       AdPlay
Description: musikseplare f�r flera format som anv�nder OPL2/3-ljud
Keywords:    adplay,adplug
End
