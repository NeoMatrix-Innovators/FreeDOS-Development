Begin3
Language:    SV, 850
Title:       DOSUTIL
Description: En samling sm� verktyg f�r kommandofiler
Keywords:    DOSUTILS SCRDUMP
End
