Begin3
Language:    SV, 850
Title:       CPI (Code Page Information)-paket
Description: Paket DISPLAY-typ, UPX-komprimerade CPI-filer f�r diverse DOS-kodsidor.
Keywords:    visa, kodsida, cp, dos kodsida, dos cp, teckenupps�ttning
End
