Begin3
Language:    SV, 850
Title:       WATTCP
Description: WATTCP
Keywords:    freedos, curl
End
