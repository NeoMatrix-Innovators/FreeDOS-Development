Begin3
Language:    SV, 850
Title:       cdrcache
Description: CD-ROM-cache, cachar l�sningar f�r en enhet, XMS, 386 eller b�ttre
Keywords:    cache, freedos, smartdrv, cd-rom
End
