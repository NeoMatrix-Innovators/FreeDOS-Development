Begin3
Language:    SV, 850
Title:       Zerofill
Description: Fyller tomt utrymme p� en enhet med nollor.
Summary:     Fyller tomt utrymme p� en enhet med nollor. Det hj�lper virtuella maskiner och programvara f�r diskkompression att komprimera allokerat utrymme p� volymen och reducerar d�rf�r dess diskanv�ndning.
Keywords:    dos
End
