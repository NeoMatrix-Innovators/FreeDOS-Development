Begin3
Language:    SV, 850
Title:       MD5SUM
Description: Ber�knar MD5 kontrollsummor
Keywords:    md5, md5sum, kontrollsumma, kryptografisk, sha, crc
End
