FD-REPOv1	Build time: 1645361091	Enhetsdrivrutiner	16
cdrcache	2004-05-13a	CD-ROM-cache, cachar l�sningar f�r en enhet, XMS, 386 eller b�ttre	2484bd2a
doslfn	0.41d	Tillhandah�ller LFN (L�nga FilNamn) API:et i ren DOS (utan Windows)	8726041d
gcdrom	2.4b	SATA inbyggd IDE CD/DVD-ROM-drivrutin f�r DOS (ocks� k�nd som 'ODD DOS-drivrutin') med st�d f�r alla SATA inbyggda IDE-styrkort s� som Intel ICH6/ICH7/ICH8, Jmicron 363/368, Nvidia CK804 MCP55/MCP51 etc. (byggt fr�n XCDROM med �ndrat namn)	63fb5de0
hiram	1.9a	�vre minnesut�kare (UMB) f�r 80286, 80386, 80486 CPU:er	550728b5
lfndos	1.06a	Tillhandah�ller Windows 95:s API f�r l�nga filnamn till DOS-program. DOS-program som kan anv�nda l�nga filnamn, till exempel DOS 7 Command.com, edit.com och alla DJGPP-program kan l�sa in och spara dem med hj�lp av LFNDOS. Designat f�r Win95-anv�ndare som anv�nder DOS-l�ge, men det fungerar �ven under �ldre DOS-versioner.	2a0a4419
lptdrv	0.7a	Ett verktyg f�r att styra LPT-anslutna enheter manuellt eller p� tidsbasis	50863821
ntfs	30Mar2001 (rev A)	M�jligg�r �tkomst av NTFS-partitioner	362ef6db
shareext	2.0a	Share Extender	d4f54b79
shsufdrv	1.02a	SHSUFDRV �r en drivrutin f�r diskett- och h�rddiskavbildningar. SHSURDRV kopierar avbildningen till RAM och/eller skapar RAM-enheter.	d62292b1
spool	2.2a	Spolar filutskrifter i bakgrunden. Detta kr�ver inte anv�ndning av PRINT-kommandot.	9597704c
srdisk	2.09d	Ramdisk som kan �ndra storlek. Srdisk �r en snabb och kan anv�nd mer �n 32MB XMS och EMS-minne. Storleken p� disket kan �ndras utan att starta och eller att f�rlora inneh�ll. Kompatibel med diskcopy.	db1a819e
udvd2	2015-03-05d	CD/DVD UltraDMA-enhetsdrivrutin	f17eefb5
uhdd	2021-10-30	UHDD �r en cachande drivrutin f�r upp till 10 BIOS h�rddiskar/SSD p� upp till 4 UltraDMA-styrkort. Det kommer ocks� att tillhandah�lla cachning f�r diskar som hanteras av UDVD2 om det l�ses in efter UHDD.	18c6e633
uide	2020-07-07a	En cachande drivrutin f�r allm�nt bruk f�r DOS-enheter, diskett, CD/DVD, SATA och UltraDMA-diskar	8ce0e4b3
usbdos	2010-01-30a	Samling DOS-drivrutiner f�r UHCI (USB 1.1 12Mbit/1.5Mbit)	47a59627
xkeyb	1.15a	Tangentbordsdrivrutin f�r internationellt st�d. Inkluderar ocks� KEYMAN + KLIB + LISTXDEF + SCANKBD	c1e50ea2
