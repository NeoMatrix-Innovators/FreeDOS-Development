Begin3
Language:    SV, 850
Title:       setedit
Description: En textredigerare f�r programmerare f�r DJGPP, liknar BC++ IDE och RHIDE
Summary:     setedit �r en v�nlig textredigerare f�r konsolen med utseende och k�nsla fr�n Borlands redigerare f�r DOS. Denna manualsidal beskriver endast kommandoradsflaggorna f�r redigeraren. Du kan f�r fullst�ndig hj�lp om redigeraren genom att anv�nda hj�lpen i redigeraren. Ett godtyckligt antal filnamn kan komma efter flaggorna och de kommer automatiskt att l�sas in av redigeraren i samma ordning som du anger dem. Du kan ange extra kommandoradsflaggor via milj�variabeln SET_CMD-LINE. L�s dokumentation f�r vidare information om denna funktion. (Notera: setedit kan inte k�ra under DOSBox)
Keywords:    redigerare, unicode, DJGPP
End
