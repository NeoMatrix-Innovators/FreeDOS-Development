Begin3
Language:    SV, 850
Title:       e3
Description: En liten textredigerarer som finns i b�de 32- och 16-bitars versioner
Keywords:    redigerare
End
