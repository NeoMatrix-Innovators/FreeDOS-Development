Begin3
Language:    SV, 850
Title:       b64
Description: Verktyg som implementerat Content-Transfer-Encoding-standarden Base64 beskriven i RFC1113.
Keywords:    b64,base64
End
