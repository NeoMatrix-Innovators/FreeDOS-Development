Begin3
Language:    SV, 850
Title:       localcfg
Description: Konfigurationsverktyg f�r lokalinst�llningar
Keywords:    country.sys
End
