Begin3
Language:    SV, 850
Title:       SHARE
Description: Installerar fildelning och l�sningsm�jligheter p� din h�rddisk - endast f�r FreeDOS-k�rnan
Keywords:    delning,fildelning
End
