Begin3
Language:    SV, 850
Title:       xDel
Description: Ut�kad filborttagning, liknar DR-DOS
Keywords:    xdel, del, deltree, ta bort
End
