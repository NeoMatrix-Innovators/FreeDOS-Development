Begin3
Language:    SV, 850
Title:       GNU sed
Description: GNU sed �r en GNU-implementation av POSIX str�mredigerarer `sed'.
Keywords:    sed
End
