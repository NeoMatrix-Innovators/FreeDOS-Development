Begin3
Language:    SV, 850
Title:       MSKERMIT
Description: Kommunikationssvit fr�n Columbia universitetet.
Summary:     MS-DOS Kermit programvarupaket f�r kommunikation f�r IBM PC och kompatibler erbjuder en upps�ttning terminalemuleringar, seriella och n�tverksbaserade kommunikationsmetoder internationell teckenkonvertering, skriptningssp�rk och Kermit fil�verf�ring.
Keywords:    serie,kommunikation,terminal,fil�verf�ring
End
