Begin3
Language:    SV, 850
Title:       DOS Navigator 2
Description: DOS Navigator 2 �ppen k�llkod�r en filhanterare baserad p� DOS Navigator (c) 1991-99 av RIT Research Labs.
Keywords:    dos navigator, norton commander
End
