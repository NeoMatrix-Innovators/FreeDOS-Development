Begin3
Language:    SV, 850
Title:       Nasm
Description: Netwide Assembler (UPX-komprimerad version)
Summary:     Netwide Assembler, NASM, �r en 80x86 och x86-64 assemblator designad f�r portabilitet och modularitet. Den har st�d f�r en uppsj� objektfilsformat, inklusive Linux och *BSD a.out, ELF, COFF, Mach-O, 16- och 32-bitars OBJ (OMF) format, Win32 och Win64. Den kan ocks� mata ut rena bin�rfiler, Intel hex- och Motorola S-Record-format. Dess syntax �r designad f�r att vara enkel och l�tt att f�rst�, likna syntaxen i Intels programutvecklingsmanual med minimal complexitet. Den har st�d f�r alla k�nda x86-arkitekturtill�gg och har bra st�d f�r makron.
Keywords:    nasm, asm, assemblator, assembler
End
