Begin3
Language:    SV, 850
Title:       SLOWDOWN
Description: G�r en snabb dator l�ngsammare. Hastigheten �r helt konfigurerbar fr�n kommandoraden eller med hj�lp av snabbtangenter. Har flera olika s�tt eller l�gen f�r att g�ra datorn l�ngsammare.
Keywords:    DOS
End
