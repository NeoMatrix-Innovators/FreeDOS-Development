Begin3
Language:    SV, 850
Title:       LBACACHE
Description: Diskcache, cachar l�sningar f�r upp till 8 CHS/LBA-h�rddiskar och disketter. XMS, 386 eller b�ttre - lbacache f�ljer med tickle!
Keywords:    cache, smartdrv, nwcache
End
