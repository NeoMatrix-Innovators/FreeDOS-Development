Begin3
Language:    SV, 850
Title:       UnRTF
Description: Konverterar dokument i RTF-format till andra format (html,latex,txt...)
Keywords:    rtf
End
