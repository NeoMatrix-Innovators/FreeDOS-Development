Begin3
Language:    SV, 850
Title:       GZIP
Description: GNU zip-komprimering - ett filarkvieringsverktyg, i stil med PKZIP
Keywords:    gzip, zip, unzip, arkivprogram, packer
End
