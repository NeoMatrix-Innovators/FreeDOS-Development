Begin3
Language:    SV, 850
Title:       MinEd
Description: Textredigerare med utf�rligt Unicode- och CJK-st�d. Beh�ndig och effktiva funktioner f�r redigering av rena textdokument, program, HTML, osv. Anv�ndarv�ndligt gr�nssnitt, musstyrning och menyer.
Summary:     Mined �r en kraftfull textredigerare. Mined tillhandah�ller b�de omfattande Unicode- och CJK-st�d med st�d f�r m�nga specifika funktioner och t�cker specialfall som �ndra redigerare inte �r medvetna om (s� som autoidetifieringsfunktion och automatiskt hantering av terminalvarianter eller Han-tecken information). Det var den f�rsta redigeraren som hade st�d f�r Unicode i en ren textterminal (som xterm eller rxvt).
Keywords:    redigera, redigerare, unicode, kodsida, kodning
End
