Begin3
Language:    SV, 850
Title:       CWSDPMI
Description: 32-bitars DPI DOS extender designad f�r DJGPP.
Keywords:    extender, DPMI, DJGPP
End
