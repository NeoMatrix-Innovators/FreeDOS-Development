Begin3
Language:    SV, 850
Title:       BSUM
Description: ber�knar BSD-kontrollsummor f�r filer
Summary:     bsum �r ett litet verktyg (256 byte!) som ber�knar BSD-kontrollsummor
Keywords:    dos
End
