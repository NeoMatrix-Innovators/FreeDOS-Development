Begin3
Language:    SV, 850
Title:       bmp2png
Description: Kommandoradsverktyg som konverterar BMP-bilder till PNG (och omv�nt)
Keywords:    bmp,png
End
